2,26483
712
83
0
0
0
4
5
0
0
0
0,09
1,48
2
6
10
0,44
0,3
0,66
3
1
1,35
True
True
False
False
False
